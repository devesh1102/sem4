library std;
use std.textio.all;
 
library std;
use std.standard.all;
 
library ieee;
use ieee.std_logic_1164.all;
 
entity Testbench is
end entity;
architecture Behave of Testbench is
 
  ----------------------------------------------------------------
  --  edit the following lines to set the number of i/o's of your
  --  DUT.
  ----------------------------------------------------------------
  constant number_of_inputs  : integer := 7;  -- # input bits to your design.
  constant number_of_outputs : integer := 1;  -- # output bits from your design.
 
  -- component port widths..
  component DUT is
   port(input_vector: in std_logic_vector(number_of_inputs-1  downto 0);   
        output_vector: out std_logic_vector(number_of_outputs-1 downto 0));
  end component;
 
  -- end editing.
  ----------------------------------------------------------------
  ----------------------------------------------------------------
 
  signal input_vector  : std_logic_vector(number_of_inputs-1 downto 0);
  signal output_vector : std_logic_vector(number_of_outputs-1 downto 0);
 
  -- create a constrained string outof
  function to_string(x: string) return string is
      variable ret_val: string(1 to x'length);
      alias lx : string (1 to x'length) is x;
  begin 
      ret_val := lx;
      return(ret_val);
  end to_string;
 
begin
  process
    variable err_flag : boolean := false;
	 ----------------------------------------------------------------------------
	 --add address of tracefile and output 
    File INFILE: text open read_mode is "/home/student/devesh/string_new/string_recognizer_test_files/tracefile1.txt";
    FILE OUTFILE: text  open write_mode is "/home/student/devesh/string_new/string_recognizer_test_files/OUTPUT1pc1.txt";
 
    ---------------------------------------------------
    -- edit the next two lines to customize
    ---------------------------------------------------
    variable input_vector_var: bit_vector (number_of_inputs-1 downto 0);
    variable output_vector_var: bit_vector (number_of_outputs-1 downto 0);
    variable output_mask_var: bit_vector (number_of_outputs-1 downto 0);
    variable output_comp_var: bit_vector (number_of_outputs-1 downto 0);
    constant ZZZZ : bit_vector(number_of_outputs-1 downto 0) := (others => '0');
    ----------------------------------------------------
 
    variable INPUT_LINE: Line;
    variable OUTPUT_LINE: Line;
    variable LINE_COUNT: integer := 0;
 
   
  begin
    while not endfile(INFILE) loop
          -- will read a new line every 5ns, apply input,
          -- wait for 1 ns for circuit to settle.
          -- read output.
 
 
          LINE_COUNT := LINE_COUNT + 1;
 
 
          -- read input at current time.
          readLine (INFILE, INPUT_LINE);
          read (INPUT_LINE, input_vector_var);
          read (INPUT_LINE, output_vector_var);
          read (INPUT_LINE, output_mask_var);
       
          -- apply input.
          input_vector <= to_stdlogicvector(input_vector_var);
 
          -- wait for the circuit to settle
          wait for 1 ns;
 
          -- check output.
          output_comp_var := (output_mask_var and (to_bitvector(output_vector) xor output_vector_var));
          if (output_comp_var  /= ZZZZ) then
             write(OUTPUT_LINE,to_string("ERROR: line "));
             write(OUTPUT_LINE, LINE_COUNT);
             writeline(OUTFILE, OUTPUT_LINE);
             err_flag := true;
          end if;
 
          write(OUTPUT_LINE, to_bitvector(input_vector));
          write(OUTPUT_LINE, to_string(" "));
          write(OUTPUT_LINE, to_bitvector(output_vector));
          writeline(OUTFILE, OUTPUT_LINE);
 
          -- advance time by 4 ns.
          wait for 1 ns;
    end loop;
 
    assert (err_flag) report "SUCCESS, all tests passed." severity note;
    assert (not err_flag) report "FAILURE, some tests failed." severity error;
 
    wait;
  end process;
 
  dut_instance: DUT
        port map(input_vector => input_vector, output_vector =>output_vector );
 
end Behave;
